
// Group N0.- 09
//Group name - Inteljr
//LAB - 3 - Memory block for microprocessor 
//date - 1/09/16

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:05:59 09/04/2016 
// Design Name: 
// Module Name:    Data_mem 
// Project Name: 	Data memory block for microprocessor 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Data_mem(mux_ans_dm,RW_dm,ans_ex,B_Bypass,RW_ex,mem_en_ex,mem_rw_ex,mem_mux_sel_ex,clk,reset );

//outputs
output [7:0]mux_ans_dm;
output reg [4:0]RW_dm;
//inputs
input [7:0]ans_ex,B_Bypass;
input [4:0]RW_ex;
input  mem_en_ex,mem_rw_ex,mem_mux_sel_ex,clk,reset;

reg mem_mux_sel_dm;
reg [7:0]ans_reg;
wire [4:0] RW_dm_temp;
wire [7:0] ans_reg_temp;
wire mem_mux_sel_dm_temp;
wire [7:0]ans_dm;

//Resetting all ouputs of data memory block 
assign RW_dm_temp = (reset==1'b1) ? RW_ex : 5'b0;
assign ans_reg_temp = (reset==1'b1) ? ans_ex : 8'b0;
assign mem_mux_sel_dm_temp = (reset==1'b1) ? mem_mux_sel_ex: 1'b0;

//Sequantial Logic
always@(posedge clk)    //Generate new instruction at every Positive Edge of clock!! 
begin 
	RW_dm <= RW_dm_temp;
	ans_reg <= ans_reg_temp;
	mem_mux_sel_dm<=mem_mux_sel_dm_temp;
end

//Instance of data memory block generated by IP core generator

DM_IM dm(
  .clka(clk), // input clka
  .ena(mem_en_ex), // input ena
  .wea(mem_rw_ex), // input [0 : 0] wea
  .addra(ans_ex), // input [7 : 0] addra
  .dina(B_Bypass), // input [7 : 0] dina
  .douta(ans_dm) // output [7 : 0] douta
);
//Combinational Logic
assign mux_ans_dm = (mem_mux_sel_dm == 1) ? ans_dm: ans_reg;//mux to select between output from register or output from data memory
endmodule


